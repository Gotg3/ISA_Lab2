library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;



package dadda_package is
    
	constant k: integer:=32;    --operand bits
	constant k_row:  integer:=33;	 --bits in the row k+1 bits
	
end package dadda_package;